library IEEE; library WORK;
use work.jpeg_Package.all;
use ieee.numeric_std.all;
entity tb is
end tb;
architecture simul of tb is
    signal quantizer_res : integer_MCU;
    signal input, fourier_res : real_MCU;
    signal zigzag_res : integer_array;
begin   
    input (0,0) <= real(-76);
    input (0,1) <= real(-73);
    input (0,2) <= real(-67);
    input (0,3) <= real(-62);
    input (0,4) <= real(-58);
    input (0,5) <= real(-67);
    input (0,6) <= real(-64);
    input (0,7) <= real(-55);
    input (1,0) <= real(-65);
    input (1,1) <= real(-69);
    input (1,2) <= real(-73);
    input (1,3) <= real(-38);
    input (1,4) <= real(-19);
    input (1,5) <= real(-43);
    input (1,6) <= real(-59);
    input (1,7) <= real(-56);
    input (2,0) <= real(-66);
    input (2,1) <= real(-69);
    input (2,2) <= real(-60);
    input (2,3) <= real(-15);
    input (2,4) <= real(16);
    input (2,5) <= real(-24);
    input (2,6) <= real(-62);
    input (2,7) <= real(-55);
    input (3,0) <= real(-65);
    input (3,1) <= real(-70);
    input (3,2) <= real(-57);
    input (3,3) <= real(-6);
    input (3,4) <= real(26);
    input (3,5) <= real(-22);
    input (3,6) <= real(-58);
    input (3,7) <= real(-59);
    input (4,0) <= real(-61);
    input (4,1) <= real(-67);
    input (4,2) <= real(-60);
    input (4,3) <= real(-24);
    input (4,4) <= real(-2);
    input (4,5) <= real(-40);
    input (4,6) <= real(-60);
    input (4,7) <= real(-58);
    input (5,0) <= real(-49);
    input (5,1) <= real(-63);
    input (5,2) <= real(-68);
    input (5,3) <= real(-58);
    input (5,4) <= real(-51);
    input (5,5) <= real(-60);
    input (5,6) <= real(-70);
    input (5,7) <= real(-53);
    input (6,0) <= real(-43);
    input (6,1) <= real(-57);
    input (6,2) <= real(-64);
    input (6,3) <= real(-69);
    input (6,4) <= real(-73);
    input (6,5) <= real(-67);
    input (6,6) <= real(-63);
    input (6,7) <= real(-45);
    input (7,0) <= real(-41);
    input (7,1) <= real(-49);
    input (7,2) <= real(-59);
    input (7,3) <= real(-60);
    input (7,4) <= real(-63);
    input (7,5) <= real(-52);
    input (7,6) <= real(-50);
    input (7,7) <= real(-34);
    process begin
        wait for 5 ns;
        fourier_res <= Fourier(input);
	    wait for 5 ns;
        quantizer_res <= Quantizer (fourier_res, Y_Quantizer_Matrix);
        wait for 5 ns;
        zigzag_res <= Zigzag(quantizer_res);
        wait;
    end process; 
end simul ;     